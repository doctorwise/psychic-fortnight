../../../mode/hdl/vhdl/mode.vhd