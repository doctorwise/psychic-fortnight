module inv(input logic a,
	   output logic y);

   assign y = ~a;

endmodule
