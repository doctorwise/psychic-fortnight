../../../4_15_structural_mux2/hdl/sv/tristate.sv