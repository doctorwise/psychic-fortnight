../../../4_15_structural_mux2/hdl/vhdl/tristate.vhd