.PHONY: all

all:
	@./.build_sv.sh
