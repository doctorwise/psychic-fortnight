../../../4_05_multiplexer/hdl/vhdl/mux2.hdl