../../../4_05_multiplexer/hdl/sv/mux2.sv