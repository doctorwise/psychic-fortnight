module and8 (
		input	logic[7:0] a,
		output	logic	   b
	);

	assign y = &a;

endmodule
