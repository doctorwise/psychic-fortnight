../../../4_15_structural_mux2/hdl/vhdl/mux2.vhd