../../../4_34_parameterizedmux2/hdl/sv/mux2.sv