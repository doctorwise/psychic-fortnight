../../../4_10_tristate/hdl/vhdl/tristate.hdl