../../../lights/hdl/sv/lights.sv