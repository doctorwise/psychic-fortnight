../../../4_34_parameterizedmux2/hdl/vhdl/mux2.vhd