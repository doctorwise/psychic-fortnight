../../../4_26_priority/hdl/vhdl/priority.vhd