../../../lights/hdl/vhdl/lights.vhd