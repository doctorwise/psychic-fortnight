../../../4_10_tristate/hdl/sv/tristate.sv