../../../mode/hdl/sv/mode.sv